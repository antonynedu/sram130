.lib "/home/antony/tools/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice" tt


XM2 Qb Q gnd! gnd! sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 m=1
XM4 Q Qb gnd! gnd! sky130_fd_pr__nfet_01v8 L=0.15 W=0.6 m=1
XM5 Q WL BL gnd! sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 m=1
XM6 Qb WL BLb gnd! sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 m=1
XM1 Qb Q vdd! vdd! sky130_fd_pr__pfet_01v8 L=0.15 W=0.3 m=1
XM3 Q Qb vdd! vdd! sky130_fd_pr__pfet_01v8 L=0.15 W=0.3 m=1


*Test Pulses
v1 BL 0 pulse(0 1.8 0ns 60ps 60ps 5ns 10ns)
v2 WL 0 dc 1.8v


**************
.tran 1e-09 20e-09 0e-00
.control
run
plot WL BL-2 BLb-4 Q-6 Qb-8


.end
